/* filename
 *
 * Copyright: Victor Wen, vic7tor@gmail.com
 * This code publish under GNU GPL License
 *
 * i2d ex module
 */

`include "i2d_defines.v"

module i2d_ex(
	rst, clk,
	//input
	id_ins, id_pc, ex_dis,
	//ouput
	mau_op, sel_mau_addr
);


endmodule

